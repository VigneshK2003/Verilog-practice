module or_gate(input a ,input b ,output y );
  or(y,a,b);
endmodule

